VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_pong
  CLASS BLOCK ;
  FOREIGN wrapped_pong ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.250 296.000 25.810 300.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 0.420 300.000 1.620 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 79.300 300.000 80.500 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 86.780 300.000 87.980 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 94.940 300.000 96.140 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 102.420 300.000 103.620 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 110.580 300.000 111.780 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 118.740 300.000 119.940 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 126.220 300.000 127.420 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 134.380 300.000 135.580 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 141.860 300.000 143.060 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 150.020 300.000 151.220 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 7.900 300.000 9.100 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 158.180 300.000 159.380 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 165.660 300.000 166.860 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 173.820 300.000 175.020 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 181.300 300.000 182.500 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 189.460 300.000 190.660 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 197.620 300.000 198.820 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.100 300.000 206.300 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 213.260 300.000 214.460 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 220.740 300.000 221.940 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 228.900 300.000 230.100 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.060 300.000 17.260 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 237.060 300.000 238.260 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.540 300.000 245.740 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 252.700 300.000 253.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 260.180 300.000 261.380 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.340 300.000 269.540 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 276.500 300.000 277.700 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 283.980 300.000 285.180 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 292.140 300.000 293.340 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.540 300.000 24.740 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 31.700 300.000 32.900 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 39.860 300.000 41.060 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 47.340 300.000 48.540 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 55.500 300.000 56.700 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 62.980 300.000 64.180 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 71.140 300.000 72.340 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 5.180 300.000 6.380 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 84.060 300.000 85.260 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 92.220 300.000 93.420 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 100.380 300.000 101.580 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.860 300.000 109.060 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 116.020 300.000 117.220 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 123.500 300.000 124.700 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 131.660 300.000 132.860 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 139.820 300.000 141.020 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 147.300 300.000 148.500 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 155.460 300.000 156.660 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 13.340 300.000 14.540 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 162.940 300.000 164.140 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 171.100 300.000 172.300 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.260 300.000 180.460 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 186.740 300.000 187.940 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 194.900 300.000 196.100 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 202.380 300.000 203.580 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 210.540 300.000 211.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 218.700 300.000 219.900 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 226.180 300.000 227.380 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 234.340 300.000 235.540 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 20.820 300.000 22.020 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 241.820 300.000 243.020 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 249.980 300.000 251.180 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.140 300.000 259.340 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 265.620 300.000 266.820 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 273.780 300.000 274.980 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 281.260 300.000 282.460 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.420 300.000 290.620 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 297.580 300.000 298.780 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 28.980 300.000 30.180 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 37.140 300.000 38.340 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.620 300.000 45.820 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 52.780 300.000 53.980 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 60.260 300.000 61.460 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 68.420 300.000 69.620 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 76.580 300.000 77.780 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 2.460 300.000 3.660 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 81.340 300.000 82.540 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 89.500 300.000 90.700 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 97.660 300.000 98.860 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 105.140 300.000 106.340 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 113.300 300.000 114.500 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 120.780 300.000 121.980 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 128.940 300.000 130.140 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 137.100 300.000 138.300 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 144.580 300.000 145.780 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 152.740 300.000 153.940 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.620 300.000 11.820 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 160.220 300.000 161.420 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 168.380 300.000 169.580 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 176.540 300.000 177.740 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 184.020 300.000 185.220 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 192.180 300.000 193.380 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 200.340 300.000 201.540 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 207.820 300.000 209.020 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 215.980 300.000 217.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 223.460 300.000 224.660 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 231.620 300.000 232.820 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 18.780 300.000 19.980 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 239.780 300.000 240.980 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 247.260 300.000 248.460 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 255.420 300.000 256.620 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 262.900 300.000 264.100 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 271.060 300.000 272.260 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 279.220 300.000 280.420 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 286.700 300.000 287.900 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 294.860 300.000 296.060 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 26.260 300.000 27.460 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 34.420 300.000 35.620 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 41.900 300.000 43.100 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 50.060 300.000 51.260 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 58.220 300.000 59.420 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.700 300.000 66.900 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.860 300.000 75.060 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.780 4.000 2.980 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.860 4.000 7.060 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.620 4.000 11.820 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.250 0.000 2.810 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 0.000 49.270 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.770 0.000 54.330 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.370 0.000 58.930 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.970 0.000 63.530 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 0.000 68.130 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.170 0.000 72.730 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 0.000 77.790 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.830 0.000 82.390 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.430 0.000 86.990 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 0.000 91.590 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.850 0.000 7.410 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.630 0.000 96.190 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.230 0.000 100.790 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.290 0.000 105.850 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.890 0.000 110.450 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.490 0.000 115.050 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 0.000 119.650 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.690 0.000 124.250 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 0.000 129.310 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 0.000 133.910 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.950 0.000 138.510 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.450 0.000 12.010 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.550 0.000 143.110 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.150 0.000 147.710 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 0.000 16.610 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.650 0.000 21.210 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.250 0.000 25.810 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.310 0.000 30.870 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.910 0.000 35.470 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.510 0.000 40.070 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 0.000 44.670 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.210 0.000 152.770 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 0.000 199.230 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.730 0.000 204.290 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.330 0.000 208.890 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.930 0.000 213.490 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.530 0.000 218.090 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.130 0.000 222.690 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 0.000 227.750 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.790 0.000 232.350 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.390 0.000 236.950 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.990 0.000 241.550 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.810 0.000 157.370 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.590 0.000 246.150 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.190 0.000 250.750 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.250 0.000 255.810 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.850 0.000 260.410 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.450 0.000 265.010 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.050 0.000 269.610 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.650 0.000 274.210 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.710 0.000 279.270 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.310 0.000 283.870 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 0.000 288.470 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.410 0.000 161.970 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.510 0.000 293.070 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.110 0.000 297.670 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.010 0.000 166.570 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 0.000 171.170 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.210 0.000 175.770 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.270 0.000 180.830 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.870 0.000 185.430 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.470 0.000 190.030 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.070 0.000 194.630 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.180 4.000 159.380 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.060 4.000 204.260 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.140 4.000 208.340 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.900 4.000 213.100 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.980 4.000 217.180 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.740 4.000 221.940 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.500 4.000 226.700 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.580 4.000 230.780 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.340 4.000 235.540 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.420 4.000 239.620 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.180 4.000 244.380 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.260 4.000 163.460 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.940 4.000 249.140 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.020 4.000 253.220 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.780 4.000 257.980 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.860 4.000 262.060 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.620 4.000 266.820 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.700 4.000 270.900 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.460 4.000 275.660 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.220 4.000 280.420 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.300 4.000 284.500 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.060 4.000 289.260 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.020 4.000 168.220 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.140 4.000 293.340 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.900 4.000 298.100 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.780 4.000 172.980 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.860 4.000 177.060 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.620 4.000 181.820 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.700 4.000 185.900 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.460 4.000 190.660 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.220 4.000 195.420 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.300 4.000 199.500 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.390 296.000 29.950 300.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.790 296.000 2.350 300.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.470 296.000 6.030 300.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.110 296.000 21.670 300.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 296.000 49.270 300.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.270 296.000 88.830 300.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.410 296.000 92.970 300.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.090 296.000 96.650 300.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.230 296.000 100.790 300.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.370 296.000 104.930 300.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.050 296.000 108.610 300.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.190 296.000 112.750 300.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 296.000 116.430 300.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.010 296.000 120.570 300.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.690 296.000 124.250 300.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.850 296.000 53.410 300.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.830 296.000 128.390 300.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 296.000 132.530 300.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.650 296.000 136.210 300.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.790 296.000 140.350 300.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.470 296.000 144.030 300.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.610 296.000 148.170 300.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.750 296.000 152.310 300.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.430 296.000 155.990 300.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.570 296.000 160.130 300.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.250 296.000 163.810 300.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.990 296.000 57.550 300.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.390 296.000 167.950 300.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.070 296.000 171.630 300.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.670 296.000 61.230 300.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.810 296.000 65.370 300.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.490 296.000 69.050 300.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.630 296.000 73.190 300.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.770 296.000 77.330 300.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 296.000 81.010 300.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.590 296.000 85.150 300.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.290 296.000 13.850 300.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.210 296.000 175.770 300.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.770 296.000 215.330 300.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.450 296.000 219.010 300.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.590 296.000 223.150 300.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.730 296.000 227.290 300.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.410 296.000 230.970 300.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.550 296.000 235.110 300.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.230 296.000 238.790 300.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.370 296.000 242.930 300.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.050 296.000 246.610 300.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.190 296.000 250.750 300.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.350 296.000 179.910 300.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.330 296.000 254.890 300.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.010 296.000 258.570 300.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.150 296.000 262.710 300.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.830 296.000 266.390 300.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.970 296.000 270.530 300.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.650 296.000 274.210 300.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.790 296.000 278.350 300.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.930 296.000 282.490 300.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.610 296.000 286.170 300.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.750 296.000 290.310 300.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.030 296.000 183.590 300.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.430 296.000 293.990 300.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.570 296.000 298.130 300.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.170 296.000 187.730 300.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.850 296.000 191.410 300.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.990 296.000 195.550 300.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 296.000 199.230 300.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.810 296.000 203.370 300.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.950 296.000 207.510 300.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.630 296.000 211.190 300.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.700 4.000 15.900 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.580 4.000 60.780 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.340 4.000 65.540 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.420 4.000 69.620 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.180 4.000 74.380 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.260 4.000 78.460 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.020 4.000 83.220 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.780 4.000 87.980 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.860 4.000 92.060 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.620 4.000 96.820 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.700 4.000 100.900 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.460 4.000 20.660 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.460 4.000 105.660 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.540 4.000 109.740 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.300 4.000 114.500 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.060 4.000 119.260 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.140 4.000 123.340 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.900 4.000 128.100 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.980 4.000 132.180 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.740 4.000 136.940 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.500 4.000 141.700 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.580 4.000 145.780 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.540 4.000 24.740 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.340 4.000 150.540 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.420 4.000 154.620 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.300 4.000 29.500 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.060 4.000 34.260 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.140 4.000 38.340 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.900 4.000 43.100 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.980 4.000 47.180 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.740 4.000 51.940 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.820 4.000 56.020 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.070 296.000 33.630 300.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.210 296.000 37.770 300.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.890 296.000 41.450 300.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.030 296.000 45.590 300.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.610 296.000 10.170 300.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.430 296.000 17.990 300.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 297.015 288.405 ;
      LAYER met1 ;
        RECT 1.910 4.460 297.550 288.560 ;
      LAYER met2 ;
        RECT 2.630 295.720 5.190 298.365 ;
        RECT 6.310 295.720 9.330 298.365 ;
        RECT 10.450 295.720 13.010 298.365 ;
        RECT 14.130 295.720 17.150 298.365 ;
        RECT 18.270 295.720 20.830 298.365 ;
        RECT 21.950 295.720 24.970 298.365 ;
        RECT 26.090 295.720 29.110 298.365 ;
        RECT 30.230 295.720 32.790 298.365 ;
        RECT 33.910 295.720 36.930 298.365 ;
        RECT 38.050 295.720 40.610 298.365 ;
        RECT 41.730 295.720 44.750 298.365 ;
        RECT 45.870 295.720 48.430 298.365 ;
        RECT 49.550 295.720 52.570 298.365 ;
        RECT 53.690 295.720 56.710 298.365 ;
        RECT 57.830 295.720 60.390 298.365 ;
        RECT 61.510 295.720 64.530 298.365 ;
        RECT 65.650 295.720 68.210 298.365 ;
        RECT 69.330 295.720 72.350 298.365 ;
        RECT 73.470 295.720 76.490 298.365 ;
        RECT 77.610 295.720 80.170 298.365 ;
        RECT 81.290 295.720 84.310 298.365 ;
        RECT 85.430 295.720 87.990 298.365 ;
        RECT 89.110 295.720 92.130 298.365 ;
        RECT 93.250 295.720 95.810 298.365 ;
        RECT 96.930 295.720 99.950 298.365 ;
        RECT 101.070 295.720 104.090 298.365 ;
        RECT 105.210 295.720 107.770 298.365 ;
        RECT 108.890 295.720 111.910 298.365 ;
        RECT 113.030 295.720 115.590 298.365 ;
        RECT 116.710 295.720 119.730 298.365 ;
        RECT 120.850 295.720 123.410 298.365 ;
        RECT 124.530 295.720 127.550 298.365 ;
        RECT 128.670 295.720 131.690 298.365 ;
        RECT 132.810 295.720 135.370 298.365 ;
        RECT 136.490 295.720 139.510 298.365 ;
        RECT 140.630 295.720 143.190 298.365 ;
        RECT 144.310 295.720 147.330 298.365 ;
        RECT 148.450 295.720 151.470 298.365 ;
        RECT 152.590 295.720 155.150 298.365 ;
        RECT 156.270 295.720 159.290 298.365 ;
        RECT 160.410 295.720 162.970 298.365 ;
        RECT 164.090 295.720 167.110 298.365 ;
        RECT 168.230 295.720 170.790 298.365 ;
        RECT 171.910 295.720 174.930 298.365 ;
        RECT 176.050 295.720 179.070 298.365 ;
        RECT 180.190 295.720 182.750 298.365 ;
        RECT 183.870 295.720 186.890 298.365 ;
        RECT 188.010 295.720 190.570 298.365 ;
        RECT 191.690 295.720 194.710 298.365 ;
        RECT 195.830 295.720 198.390 298.365 ;
        RECT 199.510 295.720 202.530 298.365 ;
        RECT 203.650 295.720 206.670 298.365 ;
        RECT 207.790 295.720 210.350 298.365 ;
        RECT 211.470 295.720 214.490 298.365 ;
        RECT 215.610 295.720 218.170 298.365 ;
        RECT 219.290 295.720 222.310 298.365 ;
        RECT 223.430 295.720 226.450 298.365 ;
        RECT 227.570 295.720 230.130 298.365 ;
        RECT 231.250 295.720 234.270 298.365 ;
        RECT 235.390 295.720 237.950 298.365 ;
        RECT 239.070 295.720 242.090 298.365 ;
        RECT 243.210 295.720 245.770 298.365 ;
        RECT 246.890 295.720 249.910 298.365 ;
        RECT 251.030 295.720 254.050 298.365 ;
        RECT 255.170 295.720 257.730 298.365 ;
        RECT 258.850 295.720 261.870 298.365 ;
        RECT 262.990 295.720 265.550 298.365 ;
        RECT 266.670 295.720 269.690 298.365 ;
        RECT 270.810 295.720 273.370 298.365 ;
        RECT 274.490 295.720 277.510 298.365 ;
        RECT 278.630 295.720 281.650 298.365 ;
        RECT 282.770 295.720 285.330 298.365 ;
        RECT 286.450 295.720 289.470 298.365 ;
        RECT 290.590 295.720 293.150 298.365 ;
        RECT 294.270 295.720 297.290 298.365 ;
        RECT 1.940 4.280 297.520 295.720 ;
        RECT 1.940 2.195 1.970 4.280 ;
        RECT 3.090 2.195 6.570 4.280 ;
        RECT 7.690 2.195 11.170 4.280 ;
        RECT 12.290 2.195 15.770 4.280 ;
        RECT 16.890 2.195 20.370 4.280 ;
        RECT 21.490 2.195 24.970 4.280 ;
        RECT 26.090 2.195 30.030 4.280 ;
        RECT 31.150 2.195 34.630 4.280 ;
        RECT 35.750 2.195 39.230 4.280 ;
        RECT 40.350 2.195 43.830 4.280 ;
        RECT 44.950 2.195 48.430 4.280 ;
        RECT 49.550 2.195 53.490 4.280 ;
        RECT 54.610 2.195 58.090 4.280 ;
        RECT 59.210 2.195 62.690 4.280 ;
        RECT 63.810 2.195 67.290 4.280 ;
        RECT 68.410 2.195 71.890 4.280 ;
        RECT 73.010 2.195 76.950 4.280 ;
        RECT 78.070 2.195 81.550 4.280 ;
        RECT 82.670 2.195 86.150 4.280 ;
        RECT 87.270 2.195 90.750 4.280 ;
        RECT 91.870 2.195 95.350 4.280 ;
        RECT 96.470 2.195 99.950 4.280 ;
        RECT 101.070 2.195 105.010 4.280 ;
        RECT 106.130 2.195 109.610 4.280 ;
        RECT 110.730 2.195 114.210 4.280 ;
        RECT 115.330 2.195 118.810 4.280 ;
        RECT 119.930 2.195 123.410 4.280 ;
        RECT 124.530 2.195 128.470 4.280 ;
        RECT 129.590 2.195 133.070 4.280 ;
        RECT 134.190 2.195 137.670 4.280 ;
        RECT 138.790 2.195 142.270 4.280 ;
        RECT 143.390 2.195 146.870 4.280 ;
        RECT 147.990 2.195 151.930 4.280 ;
        RECT 153.050 2.195 156.530 4.280 ;
        RECT 157.650 2.195 161.130 4.280 ;
        RECT 162.250 2.195 165.730 4.280 ;
        RECT 166.850 2.195 170.330 4.280 ;
        RECT 171.450 2.195 174.930 4.280 ;
        RECT 176.050 2.195 179.990 4.280 ;
        RECT 181.110 2.195 184.590 4.280 ;
        RECT 185.710 2.195 189.190 4.280 ;
        RECT 190.310 2.195 193.790 4.280 ;
        RECT 194.910 2.195 198.390 4.280 ;
        RECT 199.510 2.195 203.450 4.280 ;
        RECT 204.570 2.195 208.050 4.280 ;
        RECT 209.170 2.195 212.650 4.280 ;
        RECT 213.770 2.195 217.250 4.280 ;
        RECT 218.370 2.195 221.850 4.280 ;
        RECT 222.970 2.195 226.910 4.280 ;
        RECT 228.030 2.195 231.510 4.280 ;
        RECT 232.630 2.195 236.110 4.280 ;
        RECT 237.230 2.195 240.710 4.280 ;
        RECT 241.830 2.195 245.310 4.280 ;
        RECT 246.430 2.195 249.910 4.280 ;
        RECT 251.030 2.195 254.970 4.280 ;
        RECT 256.090 2.195 259.570 4.280 ;
        RECT 260.690 2.195 264.170 4.280 ;
        RECT 265.290 2.195 268.770 4.280 ;
        RECT 269.890 2.195 273.370 4.280 ;
        RECT 274.490 2.195 278.430 4.280 ;
        RECT 279.550 2.195 283.030 4.280 ;
        RECT 284.150 2.195 287.630 4.280 ;
        RECT 288.750 2.195 292.230 4.280 ;
        RECT 293.350 2.195 296.830 4.280 ;
      LAYER met3 ;
        RECT 4.400 297.180 295.600 298.345 ;
        RECT 4.400 296.500 296.000 297.180 ;
        RECT 4.000 296.460 296.000 296.500 ;
        RECT 4.000 294.460 295.600 296.460 ;
        RECT 4.000 293.740 296.000 294.460 ;
        RECT 4.400 291.740 295.600 293.740 ;
        RECT 4.000 291.020 296.000 291.740 ;
        RECT 4.000 289.660 295.600 291.020 ;
        RECT 4.400 289.020 295.600 289.660 ;
        RECT 4.400 288.300 296.000 289.020 ;
        RECT 4.400 287.660 295.600 288.300 ;
        RECT 4.000 286.300 295.600 287.660 ;
        RECT 4.000 285.580 296.000 286.300 ;
        RECT 4.000 284.900 295.600 285.580 ;
        RECT 4.400 283.580 295.600 284.900 ;
        RECT 4.400 282.900 296.000 283.580 ;
        RECT 4.000 282.860 296.000 282.900 ;
        RECT 4.000 280.860 295.600 282.860 ;
        RECT 4.000 280.820 296.000 280.860 ;
        RECT 4.400 278.820 295.600 280.820 ;
        RECT 4.000 278.100 296.000 278.820 ;
        RECT 4.000 276.100 295.600 278.100 ;
        RECT 4.000 276.060 296.000 276.100 ;
        RECT 4.400 275.380 296.000 276.060 ;
        RECT 4.400 274.060 295.600 275.380 ;
        RECT 4.000 273.380 295.600 274.060 ;
        RECT 4.000 272.660 296.000 273.380 ;
        RECT 4.000 271.300 295.600 272.660 ;
        RECT 4.400 270.660 295.600 271.300 ;
        RECT 4.400 269.940 296.000 270.660 ;
        RECT 4.400 269.300 295.600 269.940 ;
        RECT 4.000 267.940 295.600 269.300 ;
        RECT 4.000 267.220 296.000 267.940 ;
        RECT 4.400 265.220 295.600 267.220 ;
        RECT 4.000 264.500 296.000 265.220 ;
        RECT 4.000 262.500 295.600 264.500 ;
        RECT 4.000 262.460 296.000 262.500 ;
        RECT 4.400 261.780 296.000 262.460 ;
        RECT 4.400 260.460 295.600 261.780 ;
        RECT 4.000 259.780 295.600 260.460 ;
        RECT 4.000 259.740 296.000 259.780 ;
        RECT 4.000 258.380 295.600 259.740 ;
        RECT 4.400 257.740 295.600 258.380 ;
        RECT 4.400 257.020 296.000 257.740 ;
        RECT 4.400 256.380 295.600 257.020 ;
        RECT 4.000 255.020 295.600 256.380 ;
        RECT 4.000 254.300 296.000 255.020 ;
        RECT 4.000 253.620 295.600 254.300 ;
        RECT 4.400 252.300 295.600 253.620 ;
        RECT 4.400 251.620 296.000 252.300 ;
        RECT 4.000 251.580 296.000 251.620 ;
        RECT 4.000 249.580 295.600 251.580 ;
        RECT 4.000 249.540 296.000 249.580 ;
        RECT 4.400 248.860 296.000 249.540 ;
        RECT 4.400 247.540 295.600 248.860 ;
        RECT 4.000 246.860 295.600 247.540 ;
        RECT 4.000 246.140 296.000 246.860 ;
        RECT 4.000 244.780 295.600 246.140 ;
        RECT 4.400 244.140 295.600 244.780 ;
        RECT 4.400 243.420 296.000 244.140 ;
        RECT 4.400 242.780 295.600 243.420 ;
        RECT 4.000 241.420 295.600 242.780 ;
        RECT 4.000 241.380 296.000 241.420 ;
        RECT 4.000 240.020 295.600 241.380 ;
        RECT 4.400 239.380 295.600 240.020 ;
        RECT 4.400 238.660 296.000 239.380 ;
        RECT 4.400 238.020 295.600 238.660 ;
        RECT 4.000 236.660 295.600 238.020 ;
        RECT 4.000 235.940 296.000 236.660 ;
        RECT 4.400 233.940 295.600 235.940 ;
        RECT 4.000 233.220 296.000 233.940 ;
        RECT 4.000 231.220 295.600 233.220 ;
        RECT 4.000 231.180 296.000 231.220 ;
        RECT 4.400 230.500 296.000 231.180 ;
        RECT 4.400 229.180 295.600 230.500 ;
        RECT 4.000 228.500 295.600 229.180 ;
        RECT 4.000 227.780 296.000 228.500 ;
        RECT 4.000 227.100 295.600 227.780 ;
        RECT 4.400 225.780 295.600 227.100 ;
        RECT 4.400 225.100 296.000 225.780 ;
        RECT 4.000 225.060 296.000 225.100 ;
        RECT 4.000 223.060 295.600 225.060 ;
        RECT 4.000 222.340 296.000 223.060 ;
        RECT 4.400 220.340 295.600 222.340 ;
        RECT 4.000 220.300 296.000 220.340 ;
        RECT 4.000 218.300 295.600 220.300 ;
        RECT 4.000 217.580 296.000 218.300 ;
        RECT 4.400 215.580 295.600 217.580 ;
        RECT 4.000 214.860 296.000 215.580 ;
        RECT 4.000 213.500 295.600 214.860 ;
        RECT 4.400 212.860 295.600 213.500 ;
        RECT 4.400 212.140 296.000 212.860 ;
        RECT 4.400 211.500 295.600 212.140 ;
        RECT 4.000 210.140 295.600 211.500 ;
        RECT 4.000 209.420 296.000 210.140 ;
        RECT 4.000 208.740 295.600 209.420 ;
        RECT 4.400 207.420 295.600 208.740 ;
        RECT 4.400 206.740 296.000 207.420 ;
        RECT 4.000 206.700 296.000 206.740 ;
        RECT 4.000 204.700 295.600 206.700 ;
        RECT 4.000 204.660 296.000 204.700 ;
        RECT 4.400 203.980 296.000 204.660 ;
        RECT 4.400 202.660 295.600 203.980 ;
        RECT 4.000 201.980 295.600 202.660 ;
        RECT 4.000 201.940 296.000 201.980 ;
        RECT 4.000 199.940 295.600 201.940 ;
        RECT 4.000 199.900 296.000 199.940 ;
        RECT 4.400 199.220 296.000 199.900 ;
        RECT 4.400 197.900 295.600 199.220 ;
        RECT 4.000 197.220 295.600 197.900 ;
        RECT 4.000 196.500 296.000 197.220 ;
        RECT 4.000 195.820 295.600 196.500 ;
        RECT 4.400 194.500 295.600 195.820 ;
        RECT 4.400 193.820 296.000 194.500 ;
        RECT 4.000 193.780 296.000 193.820 ;
        RECT 4.000 191.780 295.600 193.780 ;
        RECT 4.000 191.060 296.000 191.780 ;
        RECT 4.400 189.060 295.600 191.060 ;
        RECT 4.000 188.340 296.000 189.060 ;
        RECT 4.000 186.340 295.600 188.340 ;
        RECT 4.000 186.300 296.000 186.340 ;
        RECT 4.400 185.620 296.000 186.300 ;
        RECT 4.400 184.300 295.600 185.620 ;
        RECT 4.000 183.620 295.600 184.300 ;
        RECT 4.000 182.900 296.000 183.620 ;
        RECT 4.000 182.220 295.600 182.900 ;
        RECT 4.400 180.900 295.600 182.220 ;
        RECT 4.400 180.860 296.000 180.900 ;
        RECT 4.400 180.220 295.600 180.860 ;
        RECT 4.000 178.860 295.600 180.220 ;
        RECT 4.000 178.140 296.000 178.860 ;
        RECT 4.000 177.460 295.600 178.140 ;
        RECT 4.400 176.140 295.600 177.460 ;
        RECT 4.400 175.460 296.000 176.140 ;
        RECT 4.000 175.420 296.000 175.460 ;
        RECT 4.000 173.420 295.600 175.420 ;
        RECT 4.000 173.380 296.000 173.420 ;
        RECT 4.400 172.700 296.000 173.380 ;
        RECT 4.400 171.380 295.600 172.700 ;
        RECT 4.000 170.700 295.600 171.380 ;
        RECT 4.000 169.980 296.000 170.700 ;
        RECT 4.000 168.620 295.600 169.980 ;
        RECT 4.400 167.980 295.600 168.620 ;
        RECT 4.400 167.260 296.000 167.980 ;
        RECT 4.400 166.620 295.600 167.260 ;
        RECT 4.000 165.260 295.600 166.620 ;
        RECT 4.000 164.540 296.000 165.260 ;
        RECT 4.000 163.860 295.600 164.540 ;
        RECT 4.400 162.540 295.600 163.860 ;
        RECT 4.400 161.860 296.000 162.540 ;
        RECT 4.000 161.820 296.000 161.860 ;
        RECT 4.000 159.820 295.600 161.820 ;
        RECT 4.000 159.780 296.000 159.820 ;
        RECT 4.400 157.780 295.600 159.780 ;
        RECT 4.000 157.060 296.000 157.780 ;
        RECT 4.000 155.060 295.600 157.060 ;
        RECT 4.000 155.020 296.000 155.060 ;
        RECT 4.400 154.340 296.000 155.020 ;
        RECT 4.400 153.020 295.600 154.340 ;
        RECT 4.000 152.340 295.600 153.020 ;
        RECT 4.000 151.620 296.000 152.340 ;
        RECT 4.000 150.940 295.600 151.620 ;
        RECT 4.400 149.620 295.600 150.940 ;
        RECT 4.400 148.940 296.000 149.620 ;
        RECT 4.000 148.900 296.000 148.940 ;
        RECT 4.000 146.900 295.600 148.900 ;
        RECT 4.000 146.180 296.000 146.900 ;
        RECT 4.400 144.180 295.600 146.180 ;
        RECT 4.000 143.460 296.000 144.180 ;
        RECT 4.000 142.100 295.600 143.460 ;
        RECT 4.400 141.460 295.600 142.100 ;
        RECT 4.400 141.420 296.000 141.460 ;
        RECT 4.400 140.100 295.600 141.420 ;
        RECT 4.000 139.420 295.600 140.100 ;
        RECT 4.000 138.700 296.000 139.420 ;
        RECT 4.000 137.340 295.600 138.700 ;
        RECT 4.400 136.700 295.600 137.340 ;
        RECT 4.400 135.980 296.000 136.700 ;
        RECT 4.400 135.340 295.600 135.980 ;
        RECT 4.000 133.980 295.600 135.340 ;
        RECT 4.000 133.260 296.000 133.980 ;
        RECT 4.000 132.580 295.600 133.260 ;
        RECT 4.400 131.260 295.600 132.580 ;
        RECT 4.400 130.580 296.000 131.260 ;
        RECT 4.000 130.540 296.000 130.580 ;
        RECT 4.000 128.540 295.600 130.540 ;
        RECT 4.000 128.500 296.000 128.540 ;
        RECT 4.400 127.820 296.000 128.500 ;
        RECT 4.400 126.500 295.600 127.820 ;
        RECT 4.000 125.820 295.600 126.500 ;
        RECT 4.000 125.100 296.000 125.820 ;
        RECT 4.000 123.740 295.600 125.100 ;
        RECT 4.400 123.100 295.600 123.740 ;
        RECT 4.400 122.380 296.000 123.100 ;
        RECT 4.400 121.740 295.600 122.380 ;
        RECT 4.000 120.380 295.600 121.740 ;
        RECT 4.000 120.340 296.000 120.380 ;
        RECT 4.000 119.660 295.600 120.340 ;
        RECT 4.400 118.340 295.600 119.660 ;
        RECT 4.400 117.660 296.000 118.340 ;
        RECT 4.000 117.620 296.000 117.660 ;
        RECT 4.000 115.620 295.600 117.620 ;
        RECT 4.000 114.900 296.000 115.620 ;
        RECT 4.400 112.900 295.600 114.900 ;
        RECT 4.000 112.180 296.000 112.900 ;
        RECT 4.000 110.180 295.600 112.180 ;
        RECT 4.000 110.140 296.000 110.180 ;
        RECT 4.400 109.460 296.000 110.140 ;
        RECT 4.400 108.140 295.600 109.460 ;
        RECT 4.000 107.460 295.600 108.140 ;
        RECT 4.000 106.740 296.000 107.460 ;
        RECT 4.000 106.060 295.600 106.740 ;
        RECT 4.400 104.740 295.600 106.060 ;
        RECT 4.400 104.060 296.000 104.740 ;
        RECT 4.000 104.020 296.000 104.060 ;
        RECT 4.000 102.020 295.600 104.020 ;
        RECT 4.000 101.980 296.000 102.020 ;
        RECT 4.000 101.300 295.600 101.980 ;
        RECT 4.400 99.980 295.600 101.300 ;
        RECT 4.400 99.300 296.000 99.980 ;
        RECT 4.000 99.260 296.000 99.300 ;
        RECT 4.000 97.260 295.600 99.260 ;
        RECT 4.000 97.220 296.000 97.260 ;
        RECT 4.400 96.540 296.000 97.220 ;
        RECT 4.400 95.220 295.600 96.540 ;
        RECT 4.000 94.540 295.600 95.220 ;
        RECT 4.000 93.820 296.000 94.540 ;
        RECT 4.000 92.460 295.600 93.820 ;
        RECT 4.400 91.820 295.600 92.460 ;
        RECT 4.400 91.100 296.000 91.820 ;
        RECT 4.400 90.460 295.600 91.100 ;
        RECT 4.000 89.100 295.600 90.460 ;
        RECT 4.000 88.380 296.000 89.100 ;
        RECT 4.400 86.380 295.600 88.380 ;
        RECT 4.000 85.660 296.000 86.380 ;
        RECT 4.000 83.660 295.600 85.660 ;
        RECT 4.000 83.620 296.000 83.660 ;
        RECT 4.400 82.940 296.000 83.620 ;
        RECT 4.400 81.620 295.600 82.940 ;
        RECT 4.000 80.940 295.600 81.620 ;
        RECT 4.000 80.900 296.000 80.940 ;
        RECT 4.000 78.900 295.600 80.900 ;
        RECT 4.000 78.860 296.000 78.900 ;
        RECT 4.400 78.180 296.000 78.860 ;
        RECT 4.400 76.860 295.600 78.180 ;
        RECT 4.000 76.180 295.600 76.860 ;
        RECT 4.000 75.460 296.000 76.180 ;
        RECT 4.000 74.780 295.600 75.460 ;
        RECT 4.400 73.460 295.600 74.780 ;
        RECT 4.400 72.780 296.000 73.460 ;
        RECT 4.000 72.740 296.000 72.780 ;
        RECT 4.000 70.740 295.600 72.740 ;
        RECT 4.000 70.020 296.000 70.740 ;
        RECT 4.400 68.020 295.600 70.020 ;
        RECT 4.000 67.300 296.000 68.020 ;
        RECT 4.000 65.940 295.600 67.300 ;
        RECT 4.400 65.300 295.600 65.940 ;
        RECT 4.400 64.580 296.000 65.300 ;
        RECT 4.400 63.940 295.600 64.580 ;
        RECT 4.000 62.580 295.600 63.940 ;
        RECT 4.000 61.860 296.000 62.580 ;
        RECT 4.000 61.180 295.600 61.860 ;
        RECT 4.400 59.860 295.600 61.180 ;
        RECT 4.400 59.820 296.000 59.860 ;
        RECT 4.400 59.180 295.600 59.820 ;
        RECT 4.000 57.820 295.600 59.180 ;
        RECT 4.000 57.100 296.000 57.820 ;
        RECT 4.000 56.420 295.600 57.100 ;
        RECT 4.400 55.100 295.600 56.420 ;
        RECT 4.400 54.420 296.000 55.100 ;
        RECT 4.000 54.380 296.000 54.420 ;
        RECT 4.000 52.380 295.600 54.380 ;
        RECT 4.000 52.340 296.000 52.380 ;
        RECT 4.400 51.660 296.000 52.340 ;
        RECT 4.400 50.340 295.600 51.660 ;
        RECT 4.000 49.660 295.600 50.340 ;
        RECT 4.000 48.940 296.000 49.660 ;
        RECT 4.000 47.580 295.600 48.940 ;
        RECT 4.400 46.940 295.600 47.580 ;
        RECT 4.400 46.220 296.000 46.940 ;
        RECT 4.400 45.580 295.600 46.220 ;
        RECT 4.000 44.220 295.600 45.580 ;
        RECT 4.000 43.500 296.000 44.220 ;
        RECT 4.400 41.500 295.600 43.500 ;
        RECT 4.000 41.460 296.000 41.500 ;
        RECT 4.000 39.460 295.600 41.460 ;
        RECT 4.000 38.740 296.000 39.460 ;
        RECT 4.400 36.740 295.600 38.740 ;
        RECT 4.000 36.020 296.000 36.740 ;
        RECT 4.000 34.660 295.600 36.020 ;
        RECT 4.400 34.020 295.600 34.660 ;
        RECT 4.400 33.300 296.000 34.020 ;
        RECT 4.400 32.660 295.600 33.300 ;
        RECT 4.000 31.300 295.600 32.660 ;
        RECT 4.000 30.580 296.000 31.300 ;
        RECT 4.000 29.900 295.600 30.580 ;
        RECT 4.400 28.580 295.600 29.900 ;
        RECT 4.400 27.900 296.000 28.580 ;
        RECT 4.000 27.860 296.000 27.900 ;
        RECT 4.000 25.860 295.600 27.860 ;
        RECT 4.000 25.140 296.000 25.860 ;
        RECT 4.400 23.140 295.600 25.140 ;
        RECT 4.000 22.420 296.000 23.140 ;
        RECT 4.000 21.060 295.600 22.420 ;
        RECT 4.400 20.420 295.600 21.060 ;
        RECT 4.400 20.380 296.000 20.420 ;
        RECT 4.400 19.060 295.600 20.380 ;
        RECT 4.000 18.380 295.600 19.060 ;
        RECT 4.000 17.660 296.000 18.380 ;
        RECT 4.000 16.300 295.600 17.660 ;
        RECT 4.400 15.660 295.600 16.300 ;
        RECT 4.400 14.940 296.000 15.660 ;
        RECT 4.400 14.300 295.600 14.940 ;
        RECT 4.000 12.940 295.600 14.300 ;
        RECT 4.000 12.220 296.000 12.940 ;
        RECT 4.400 10.220 295.600 12.220 ;
        RECT 4.000 9.500 296.000 10.220 ;
        RECT 4.000 7.500 295.600 9.500 ;
        RECT 4.000 7.460 296.000 7.500 ;
        RECT 4.400 6.780 296.000 7.460 ;
        RECT 4.400 5.460 295.600 6.780 ;
        RECT 4.000 4.780 295.600 5.460 ;
        RECT 4.000 4.060 296.000 4.780 ;
        RECT 4.000 3.380 295.600 4.060 ;
        RECT 4.400 2.215 295.600 3.380 ;
      LAYER met4 ;
        RECT 173.255 55.935 174.240 158.945 ;
        RECT 176.640 55.935 186.465 158.945 ;
  END
END wrapped_pong
END LIBRARY

